LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY cnt_n16 IS
	PORT
	(	
		CLK,CI,CLR,LOAD,UPDOWN	: IN	STD_LOGIC;
		DIN						: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		CO						: OUT	STD_LOGIC;
		Q						: OUT	STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END cnt_n16;
ARCHITECTURE a OF cnt_n16 IS
--	SIGNAL QQQ : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	
PROCESS (CLK,CLR,LOAD)
	VARIABLE QQ	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	
	IF CLR='1' 
		THEN QQ:="0000";				--OTHERS=>'0'
		ELSE IF CLK='1' AND CLK' EVENT 
				THEN IF LOAD='1' 
						THEN QQ:=DIN;	--Q<=DIN
						ELSE IF CI='1'
						THEN IF UPDOWN='1'
						THEN QQ:=QQ+1;--Q<=Q+1;QQQ<=QQQ+1;
						ELSE QQ:=QQ-1;--Q<=Q-1;
						END IF;
							--	ELSE QQ:=QQ;	
							 END IF; 		
					 END IF;
			 END IF;
  	END IF;
	Q<=QQ;			--Q<=QQQ;

IF  CI='1' --zheduan shi yinwei
		THEN IF UPDOWN='1'
				THEN IF QQ="1111"
						THEN CO<='1';
						ELSE CO<='0';
					END IF;
				ELSE IF QQ="0000"
						THEN CO<='1';
						ELSE CO<='0';
					END IF;
			END IF;
		ELSE CO<='0'; --��λ
END IF;
END PROCESS;

END a;


